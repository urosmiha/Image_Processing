module test ( testIn,testOut);

input testIn;
output wire testOut;

assign testOut = 1;

endmodule
